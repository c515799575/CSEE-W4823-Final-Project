module neural_network(pixel_in,pixel_addr,weight_memory_datain,weight_addr,result,clk,begin_sign,finish_sign,w);
input [7:0]pixel_in;
input [9:0]pixel_addr;
input [9:0]weight_memory_datain;
input [4:0]weight_addr;
input clk;
input [3:0]w;
input finish_sign,begin_sign;
output reg[3:0]result;
signal_control control_flow(finish_sign,pts_load,pts_out,weight2_rd,mac2_en,mac2_clr,bias2_rd,compare_en,clk);
input_buffer buffer(pixel_in,mac_a,finish_sign);
weight_memory memory1(weight_memory_datain,pixel_addr,weight_addr,w[0],finishi_sign,clk,data_0,data_1,data_2,data_3,data_4,data_5,data_6,data_7,data_8,data_9,data_10,data_11,data_12,data_13,data_14,data_15,data_16,data_17,data_18,data_19);
mac neu0(mac_a,data_0,neural0,clk,begin_sign,finish_sign);
mac neu1(mac_a,data_1,neural1,clk,begin_sign,finish_sign);
mac neu2(mac_a,data_2,neural2,clk,begin_sign,finish_sign);
mac neu3(mac_a,data_3,neural3,clk,begin_sign,finish_sign);
mac neu4(mac_a,data_4,neural4,clk,begin_sign,finish_sign);
mac neu5(mac_a,data_5,neural5,clk,begin_sign,finish_sign);
mac neu6(mac_a,data_6,neural6,clk,begin_sign,finish_sign);
mac neu7(mac_a,data_7,neural7,clk,begin_sign,finish_sign);
mac neu8(mac_a,data_8,neural8,clk,begin_sign,finish_sign);
mac neu9(mac_a,data_9,neural9,clk,begin_sign,finish_sign);
mac neu10(mac_a,data_10,neural10,clk,begin_sign,finish_sign);
mac neu11(mac_a,data_11,neural11,clk,begin_sign,finish_sign);
mac neu12(mac_a,data_12,neural12,clk,begin_sign,finish_sign);
mac neu13(mac_a,data_13,neural13,clk,begin_sign,finish_sign);
mac neu14(mac_a,data_14,neural14,clk,begin_sign,finish_sign);
mac neu15(mac_a,data_15,neural15,clk,begin_sign,finish_sign);
mac neu16(mac_a,data_16,neural16,clk,begin_sign,finish_sign);
mac neu17(mac_a,data_17,neural17,clk,begin_sign,finish_sign);
mac neu18(mac_a,data_18,neural18,clk,begin_sign,finish_sign);
mac neu19(mac_a,data_19,neural19,clk,begin_sign,finish_sign);
bias_memory memory2(weight_memory_datain,bias_data0,bias_data1,bias_data2,bias_data3,bias_data4,bias_data5,bias_data6,bias_data7,bias_data8,bias_data9,bias_data10,bias_data11,bias_data12,bias_data13,bias_data14,bias_data15,bias_data16,bias_data17,bias_data18,bias_data19,weight_addr,finish_sign,w[1],clk);
bias_adder bias0(neural0,bias_data0,bias_result0,clk);
bias_adder bias1(neural1,bias_data1,bias_result1,clk);
bias_adder bias2(neural2,bias_data2,bias_result2,clk);
bias_adder bias3(neural3,bias_data3,bias_result3,clk);
bias_adder bias4(neural4,bias_data4,bias_result4,clk);
bias_adder bias5(neural5,bias_data5,bias_result5,clk);
bias_adder bias6(neural6,bias_data6,bias_result6,clk);
bias_adder bias7(neural7,bias_data7,bias_result7,clk);
bias_adder bias8(neural8,bias_data8,bias_result8,clk);
bias_adder bias9(neural9,bias_data9,bias_result9,clk);
bias_adder bias10(neural0,bias_data10,bias_result10,clk);
bias_adder bias11(neural1,bias_data11,bias_result11,clk);
bias_adder bias12(neural2,bias_data12,bias_result12,clk);
bias_adder bias13(neural3,bias_data13,bias_result13,clk);
bias_adder bias14(neural4,bias_data14,bias_result14,clk);
bias_adder bias15(neural5,bias_data15,bias_result15,clk);
bias_adder bias16(neural6,bias_data16,bias_result16,clk);
bias_adder bias17(neural7,bias_data17,bias_result17,clk);
bias_adder bias18(neural8,bias_data18,bias_result18,clk);
bias_adder bias19(neural9,bias_data19,bias_result19,clk);
Relu r0(bias_result0,linear2_input0,1,clk);
Relu r1(bias_result1,linear2_input1,1,clk);
Relu r2(bias_result2,linear2_input2,1,clk);
Relu r3(bias_result3,linear2_input3,1,clk);
Relu r4(bias_result4,linear2_input4,1,clk);
Relu r5(bias_result5,linear2_input5,1,clk);
Relu r6(bias_result6,linear2_input6,1,clk);
Relu r7(bias_result7,linear2_input7,1,clk);
Relu r8(bias_result8,linear2_input8,1,clk);
Relu r9(bias_result9,linear2_input9,1,clk);
Relu r10(bias_result10,linear2_input10,1,clk);
Relu r11(bias_result11,linear2_input11,1,clk);
Relu r12(bias_result12,linear2_input12,1,clk);
Relu r13(bias_result13,linear2_input13,1,clk);
Relu r14(bias_result14,linear2_input14,1,clk);
Relu r15(bias_result15,linear2_input15,1,clk);
Relu r16(bias_result16,linear2_input16,1,clk);
Relu r17(bias_result17,linear2_input17,1,clk);
Relu r18(bias_result18,linear2_input18,1,clk);
Relu r19(bias_result19,linear2_input19,1,clk);
pts pts1(linear2_input0,linear2_input1,linear2_input2,linear2_input3,linear2_input4,linear2_input5,linear2_input6,linear2_input7,linear2_input8,linear2_input9,linear2_input10,linear2_input11,linear2_input12,linear2_input13,linear2_input14,linear2_input15,linear2_input016,linear2_input17,linear2_input18,linear2_input19,linear2,clk,pts_load,pts_out);
weight_memory_linear2 linear2_mem(weight_memory_datain,linear2_m0,linear2_m1,linear2_m2,linear2_m3,linear2_m4,linear2_m5,linear2_m6,linear2_m7,linear2_m8,linear2_m9,pixel_addr[3:0],weight_addr[3:0],weight2_rd,w[2],clk);
mac2 l2n0(linear2,linear2_m0,torelu0,clk,mac2_clr,mac2_en);
mac2 l2n1(linear2,linear2_m1,torelu1,clk,mac2_clr,mac2_en);
mac2 l2n2(linear2,linear2_m2,torelu2,clk,mac2_clr,mac2_en);
mac2 l2n3(linear2,linear2_m3,torelu3,clk,mac2_clr,mac2_en);
mac2 l2n4(linear2,linear2_m4,torelu4,clk,mac2_clr,mac2_en);
mac2 l2n5(linear2,linear2_m5,torelu5,clk,mac2_clr,mac2_en);
mac2 l2n6(linear2,linear2_m6,torelu6,clk,mac2_clr,mac2_en);
mac2 l2n7(linear2,linear2_m7,torelu7,clk,mac2_clr,mac2_en);
mac2 l2n8(linear2,linear2_m8,torelu8,clk,mac2_clr,mac2_en);
mac2 l2n9(linear2,linear2_m9,torelu9,clk,mac2_clr,mac2_en);
bias2_memory bias2_mem(weight_memory_datain,bias2_w0,bias2_w1,bias2_w2,bias2_w3,bias2_w4,bias2_w5,bias2_w6,bias2_w7,bias2_w8,bias2_w9,weight_addr[3:0],bias2_rd,w[3],clk);
bias_adder bias20(torelu0,bias2_w0,bias2_result0,clk);
bias_adder bias21(torelu1,bias2_w1,bias2_result1,clk);
bias_adder bias22(torelu2,bias2_w2,bias2_result2,clk);
bias_adder bias23(torelu3,bias2_w3,bias2_result3,clk);
bias_adder bias24(torelu4,bias2_w4,bias2_result4,clk);
bias_adder bias25(torelu5,bias2_w5,bias2_result5,clk);
bias_adder bias26(torelu6,bias2_w6,bias2_result6,clk);
bias_adder bias27(torelu7,bias2_w7,bias2_result7,clk);
bias_adder bias28(torelu8,bias2_w8,bias2_result8,clk);
bias_adder bias29(torelu9,bias2_w9,bias2_result9,clk);
Relu r20(bias2_result0,compare_input0,1,clk);
Relu r21(bias2_result1,compare_input1,1,clk);
Relu r22(bias2_result2,compare_input2,1,clk);
Relu r23(bias2_result3,compare_input3,1,clk);
Relu r24(bias2_result4,compare_input4,1,clk);
Relu r25(bias2_result5,compare_input5,1,clk);
Relu r26(bias2_result6,compare_input6,1,clk);
Relu r27(bias2_result7,compare_input7,1,clk);
Relu r28(bias2_result8,compare_input8,1,clk);
Relu r29(bias2_result9,compare_input9,1,clk);
compare(compare_input0,compare_input1,compare_input2,compare_input3,compare_input4,compare_input5,compare_input6,compare_input7,compare_input8,compare_input9,result,clk,compare_en);
endmodule
